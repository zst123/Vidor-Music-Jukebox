// Taken from https://github.com/bhagman/Tone/blob/master/Tone.h
parameter NOTE_B0  = 31;
parameter NOTE_C1  = 33;
parameter NOTE_CS1 = 35;
parameter NOTE_D1  = 37;
parameter NOTE_DS1 = 39;
parameter NOTE_E1  = 41;
parameter NOTE_F1  = 44;
parameter NOTE_FS1 = 46;
parameter NOTE_G1  = 49;
parameter NOTE_GS1 = 52;
parameter NOTE_A1  = 55;
parameter NOTE_AS1 = 58;
parameter NOTE_B1  = 62;
parameter NOTE_C2  = 65;
parameter NOTE_CS2 = 69;
parameter NOTE_D2  = 73;
parameter NOTE_DS2 = 78;
parameter NOTE_E2  = 82;
parameter NOTE_F2  = 87;
parameter NOTE_FS2 = 93;
parameter NOTE_G2  = 98;
parameter NOTE_GS2 = 104;
parameter NOTE_A2  = 110;
parameter NOTE_AS2 = 117;
parameter NOTE_B2  = 123;
parameter NOTE_C3  = 131;
parameter NOTE_CS3 = 139;
parameter NOTE_D3  = 147;
parameter NOTE_DS3 = 156;
parameter NOTE_E3  = 165;
parameter NOTE_F3  = 175;
parameter NOTE_FS3 = 185;
parameter NOTE_G3  = 196;
parameter NOTE_GS3 = 208;
parameter NOTE_A3  = 220;
parameter NOTE_AS3 = 233;
parameter NOTE_B3  = 247;
parameter NOTE_C4  = 262;
parameter NOTE_CS4 = 277;
parameter NOTE_D4  = 294;
parameter NOTE_DS4 = 311;
parameter NOTE_E4  = 330;
parameter NOTE_F4  = 349;
parameter NOTE_FS4 = 370;
parameter NOTE_G4  = 392;
parameter NOTE_GS4 = 415;
parameter NOTE_A4  = 440;
parameter NOTE_AS4 = 466;
parameter NOTE_B4  = 494;
parameter NOTE_C5  = 523;
parameter NOTE_CS5 = 554;
parameter NOTE_D5  = 587;
parameter NOTE_DS5 = 622;
parameter NOTE_E5  = 659;
parameter NOTE_F5  = 698;
parameter NOTE_FS5 = 740;
parameter NOTE_G5  = 784;
parameter NOTE_GS5 = 831;
parameter NOTE_A5  = 880;
parameter NOTE_AS5 = 932;
parameter NOTE_B5  = 988;
parameter NOTE_C6  = 1047;
parameter NOTE_CS6 = 1109;
parameter NOTE_D6  = 1175;
parameter NOTE_DS6 = 1245;
parameter NOTE_E6  = 1319;
parameter NOTE_F6  = 1397;
parameter NOTE_FS6 = 1480;
parameter NOTE_G6  = 1568;
parameter NOTE_GS6 = 1661;
parameter NOTE_A6  = 1760;
parameter NOTE_AS6 = 1865;
parameter NOTE_B6  = 1976;
parameter NOTE_C7  = 2093;
parameter NOTE_CS7 = 2217;
parameter NOTE_D7  = 2349;
parameter NOTE_DS7 = 2489;
parameter NOTE_E7  = 2637;
parameter NOTE_F7  = 2794;
parameter NOTE_FS7 = 2960;
parameter NOTE_G7  = 3136;
parameter NOTE_GS7 = 3322;
parameter NOTE_A7  = 3520;
parameter NOTE_AS7 = 3729;
parameter NOTE_B7  = 3951;
parameter NOTE_C8  = 4186;
parameter NOTE_CS8 = 4435;
parameter NOTE_D8  = 4699;
parameter NOTE_DS8 = 4978;

parameter NOTE_REST = 1;
